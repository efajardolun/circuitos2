*Circuito RLC
V1 1 0 PULSE(0 5 0 0.1us 0.1us 0.2ms 0.4ms)
RG 1 2 50
L  2 3 10m
C  3 4 1n
R  4 0 6.32455k
*R  4 0 10k
*R  4 0 1k
.end
.control
tran 0.1us 0.4ms
plot V(1) V(4)
.endc